// Top level module
module top (
    clk, reset
);
input clk, reset;


endmodule